module ROM(input [31:0] address, output [31:0] inst);

	reg [31:0] memory [255:0];

	initial begin
		memory[0] = 32'b100000_00000_00000_00000_00000000000;//-- Addi	r0	,r0	,0 -> fake command if memory 0 ignored!
		memory[1] = 32'b100000_00000_00001_00000_11000001010;//-- Addi	r1	,r0	,1546
		memory[2] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[3] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[4] = 32'b000001_00000_00001_00010_00000000000;//-- Add 	r2	,r0	,r1 
		memory[5] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[6] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[7] = 32'b000011_00000_00001_00011_00000000000;//-- sub	r3	,r0	,r1
		memory[8] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[9] = 32'b000000_00000_00000_00000_00000000000;//NOPE 
		memory[10] = 32'b000101_00010_00011_00100_00000000000;//-- And	r4	,r2	,r3	
		memory[11] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[12] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[13] = 32'b100001_00011_00101_00011_01000110100;//-- Subi	r5	,r3	,6708 
		memory[14] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[15] = 32'b000000_00000_00000_00000_00000000000;//NOPE 
		memory[16] = 32'b000110_00011_00100_00101_00000000000;//-- or	r5	,r3	,r4
		memory[17] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[18] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[19] = 32'b000111_00101_00000_00110_00000000000;//-- nor 	r6	,r5	,r0
		memory[20] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[21] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[22] = 32'b000111_00100_00000_01011_00000000000;//-- nor 	r11	,r4	,r0
		memory[23] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[24] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[25] = 32'b000011_00101_00101_00101_00000000000;//-- sub	r5	,r5	,r5 
		memory[26] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[27] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[28] = 32'b100000_00000_00001_00000_10000000000;//-- Addi 	r1	,r0	,1024    
		memory[29] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[30] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[31] = 32'b100101_00001_00010_00000_00000000000;//-- st	r2	,r1	,0      
		memory[32] = 32'b100100_00001_00101_00000_00000000000;//-- ld	r5	,r1	,0
		memory[33] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[34] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[35] = 32'b101000_00101_00000_00000_00000000011;//-- Bez	r5	,3 (it was 1)
		memory[36] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[37] = 32'b000000_00000_00000_00000_00000000000;//NOPE           
		memory[38] = 32'b001000_00101_00001_00111_00000000000;//-- xor	r7	,r5	,r1
		memory[39] = 32'b001000_00101_00001_00000_00000000000;//-- xor	r0	,r5	,r1
		memory[40] = 32'b001001_00011_01011_00111_00000000000;//-- sla	r7	,r3	,r11
		memory[41] = 32'b001010_00011_01011_01000_00000000000;//-- sll	r8	,r3	,r11
		memory[42] = 32'b001011_00011_00100_01001_00000000000;//-- sra	r9	,r3	,r4
		memory[43] = 32'b001100_00011_00100_01010_00000000000;//-- srl	r10	,r3	,r4
		memory[44] = 32'b100101_00001_00011_00000_00000000100;//-- st	r3	,r1	,4       
		memory[45] = 32'b100101_00001_00100_00000_00000001000;//-- st	r4	,r1	,8       
		memory[46] = 32'b100101_00001_00101_00000_00000001100;//-- st	r5	,r1	,12      
		memory[47] = 32'b100101_00001_00110_00000_00000010000;//-- st	r6	,r1	,16      
		memory[48] = 32'b100100_00001_01011_00000_00000000100;//-- ld	r11	,r1	,4      
		memory[49] = 32'b100101_00001_00111_00000_00000010100;//-- st	r7	,r1	,20     
		memory[50] = 32'b100101_00001_01000_00000_00000011000;//-- st	r8	,r1	,24     
		memory[51] = 32'b100101_00001_01001_00000_00000011100;//-- st	r9	,r1	,28     
		memory[52] = 32'b100101_00001_01010_00000_00000100000;//-- st	r10	,r1	,32     
		memory[53] = 32'b100101_00001_01011_00000_00000100100;//-- st	r11	,r1	,36     
		memory[54] = 32'b100000_00000_00001_00000_00000000011;//-- Addi 	r1	,r0	,3      
		memory[55] = 32'b100000_00000_00100_00000_10000000000;//-- Addi	r4	,r0	,1024   
		memory[56] = 32'b100000_00000_00010_00000_00000000000;//-- Addi 	r2	,r0	,0      
		memory[57] = 32'b100000_00000_00011_00000_00000000001;//-- Addi 	r3	,r0	,1      
		memory[58] = 32'b100000_00000_01001_00000_00000000010;//-- Addi 	r9	,r0	,2 
		memory[59] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[60] = 32'b000000_00000_00000_00000_00000000000;//NOPE    
		memory[61] = 32'b001010_00011_01001_01000_00000000000;//-- sll	r8	,r3	,r9 
		memory[62] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[63] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[64] = 32'b000001_00100_01000_01000_00000000000;//-- Add 	r8	,r4	,r8
		memory[65] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[66] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[67] = 32'b100100_01000_00101_00000_00000000000;//-- ld	r5	,r8	,0       
		memory[68] = 32'b100100_01000_00110_11111_11111111100;//-- ld	r6	,r8	,-4
		memory[69] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[70] = 32'b000000_00000_00000_00000_00000000000;//NOPE     
		memory[71] = 32'b000011_00101_00110_01001_00000000000;//-- sub 	r9	,r5	,r6 
		memory[72] = 32'b100000_00000_01010_10000_00000000000;//-- Addi 	r10	,r0	,0x8000 
		memory[73] = 32'b100000_00000_01011_00000_00000010000;//-- Addi	r11	,r0	,16 
		memory[74] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[75] = 32'b000000_00000_00000_00000_00000000000;//NOPE    
		memory[76] = 32'b001010_01010_01011_01010_00000000000;//-- sll	r10	,r1	,r11
		memory[77] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[78] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[79] = 32'b000101_01001_01010_01001_00000000000;//-- And 	r9	,r9	,r10
		memory[80] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[81] = 32'b000000_00000_00000_00000_00000000000;//NOPE 
		memory[82] = 32'b101000_01001_00000_00000_00000000100;//-- Bez	r9	,4 (it was 2) 
		memory[83] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[84] = 32'b000000_00000_00000_00000_00000000000;//NOPE        
		memory[85] = 32'b100101_01000_00101_11111_11111111100;//-- st	r5	,r8	,-4     
		memory[86] = 32'b100101_01000_00110_00000_00000000000;//-- st	r6	,r8	,0      
		memory[87] = 32'b100000_00011_00011_00000_00000000001;//-- Addi 	r3	,r3	,1 
		memory[88] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[89] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[90] = 32'b101001_00001_00011_11111_11111011111;//-- BNE	r1	,r3	,-15  -18(nope)
		memory[91] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[92] = 32'b000000_00000_00000_00000_00000000000;//NOPE  
		memory[93] = 32'b100000_00010_00010_00000_00000000001;//-- Addi r2	,r2	,1  
		memory[94] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[95] = 32'b000000_00000_00000_00000_00000000000;//NOPE    
		memory[96] = 32'b101001_00001_00010_11111_11111011000;//-- BNE	r1	,r2	,-18 -22(nope)   
		memory[97] = 32'b100000_00000_00001_00000_10000000000;//-- Addi 	r1	,r0	,1024  
		memory[98] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[99] = 32'b000000_00000_00000_00000_00000000000;//NOPE 
		memory[100] = 32'b100100_00001_00010_00000_00000000000;//-- ld	,r2	,r1	,0      
		memory[101] = 32'b100100_00001_00011_00000_00000000100;//-- ld	,r3	,r1	,4      
		memory[102] = 32'b100100_00001_00100_00000_00000001000;//-- ld	,r4	,r1	,8
		memory[103] = 32'b100100_00001_00100_00000_01000001000;//-- ld	,r4	,r1	,520 
		memory[104] = 32'b100100_00001_00100_00000_10000001000;//-- ld	,r4	,r1	,1023
		memory[105] = 32'b100100_00001_00101_00000_00000001100;//-- ld	,r5	,r1	,12     
		memory[106] = 32'b100100_00001_00110_00000_00000010000;//-- ld	,r6	,r1	,16     
		memory[107] = 32'b100100_00001_00111_00000_00000010100;//-- ld	,r7	,r1	,20     
		memory[108] = 32'b100100_00001_01000_00000_00000011000;//-- ld	,r8	,r1	,24     
		memory[109] = 32'b100100_00001_01001_00000_00000011100;//-- ld	,r9	,r1	,28     
		memory[110] = 32'b100100_00001_01010_00000_00000100000;//-- ld	,r10,r1	,32     
		memory[111] = 32'b100100_00001_01011_00000_00000100100;//-- ld	,r11,r1	,36     
		memory[112] = 32'b101010_00000_00000_11111_11111111111;//-- JMP 	-1
		memory[113] = 32'b000000_00000_00000_00000_00000000000;//NOPE
		memory[114] = 32'b000000_00000_00000_00000_00000000000;//NOPE 

	end
	assign inst = memory[address[11:2]];

endmodule